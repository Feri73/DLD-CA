module Q7_Shifter_Test();
  reg A,B,C,D,i,j,k,l;
  wire W0,W1,W3,W5,W8,W9,X0,X1,X3,X5,X8,X9,Y0,Y1,Y3,Y5,Y8,Y9,Z0,Z1,Z3,Z5,Z8,Z9;
  Q6_Shifter uut0(A,B,C,D,i,j,k,l,W0,X0,Y0,Z0);
  Q7_Shifter_1 uut1(A,B,C,D,i,j,k,l,W1,X1,Y1,Z1);
  Q7_Shifter_3 uut3(A,B,C,D,i,j,k,l,W3,X3,Y3,Z3);
  Q7_Shifter_5 uut5(A,B,C,D,i,j,k,l,W5,X5,Y5,Z5);
  wire[3:0] d;
  wire[3:0] n;
  wire[3:0] w;
  assign  d[0]=D; assign  d[1]=C; assign  d[2]=B;assign  d[3]=A;
  assign    n[0]=l;assign  n[1]=k;assign  n[2]=j;assign  n[3]=i;
  assign  W9=w[3];assign  X9=w[2];assign  Y9=w[1];assign  Z9=w[0];
  Q8_Shifter uut8(A,B,C,D,i,j,k,l,W8,X8,Y8,Z8);
  Q9_Shifter uut9(d,n,w);
  initial begin
    i=0;
    j=0;
    k=0;
    l=1;
    A=0;
    B=0;
    C=0;
    D=0;
    #100 A=1;
    #100 B=1;
    #100 C=1;
    #100 l=0;k=1;
    #100 D=1;
    #100 D=1;
    #100 j=1;k=0;
    #100 A=0;
    #100 i=1;j=0;
    #100 C=0;
    #100 i=0;j=1;
    #100 $stop;
  end
endmodule