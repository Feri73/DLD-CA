module CA2_Q11_Shifter(input[7:0] d,input[7:0] n, output[7:0] w);
  assign #(152,136) w=(n[0]?d[7:0]:(n[1]?{d[6:0],1'b0}:(n[2]?{d[5:0],2'b0}:(n[3]?{d[4:0],3'b0}:(n[4]?{d[3:0],4'b0}:(n[5]?{d[2:0],5'b0}:(n[6]?{d[1:0],6'b0}:(n[7]?{d[0:0],7'b0}:{8'b0}))))))));
endmodule