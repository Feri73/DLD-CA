module Q5_AO_Test();
  reg a,b,c;
  wire w1,w3,w5;
  Q1_AO uut1(a,b,c,w1);
  Q3_AO uut3(a,b,c,w3);
  Q5_AO uut5(a,b,c,w5);
  initial begin
    a=0;
    b=0;
    c=0;//000 w=0 delay1:17-0=17 delay3:18-0=18 delay5:13-0=13
    #30 c=1;//000->001 w=0->1 delay1:42-30=12 delay3:40-30=10 delay5:43-30=13
    #30 c=0;//001->000 w=1->0 delay1:72-60=12 delay3:70-60=10 delay5:72-60=12
    #30 b=1;//010 w=0 nochange
    #30 c=1;//010->011 w=0->1 delay1:132-120=12 delay3:130-120=10 delay5:133-120=13
    #30 c=0;//011->010 w=1->0 delay1:162-150=12 delay3:160-150=10 delay5:162-150=12
    #30 a=1;//010->110 w=0->1 delay1:199-180=19 delay3:200-180=20 delay5:198-180=18
    #30 b=0;//110->100 w=1->0 delay1:227-210=17 delay3:228-210=18 delay5:223-210=13
    #30 c=1;//100->101 w=0->1 delay1:252-240=12 delay3:250-140=10 delay5:253-140=13
    #30 c=0;//101->100 w=1->0 delay1:282-270=12 delay3:280-170=10 delay5:282-170=12
    #30 b=1;//100->110 w=0->1 delay1:319-300=19 delay3:320-300=20 delay5:317-300=17
    #30 a=0;//110->010 w=1->0 delay1:347-330=17 delay3:348-330=18 delay5:348-330=18
    #30 $stop;
  end
endmodule
