library verilog;
use verilog.vl_types.all;
entity Q3_ALU_Test is
end Q3_ALU_Test;
