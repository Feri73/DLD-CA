library verilog;
use verilog.vl_types.all;
entity Q1_Barrel_Shifter_Test is
end Q1_Barrel_Shifter_Test;
