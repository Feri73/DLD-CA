module Q2_AO_Test();
  reg a,b,c;
  wire w;
  Q1_AO uut(a,b,c,w);
  initial begin
    a=0;
    b=0;
    c=0;//000 w=0 delay:17-0=17
    #30 c=1;//000->001 w=0->1 delay:42-30=12
    #30 c=0;//001->000 w=1->0 delay:72-60=12
    #30 b=1;//010 w=0 nochange
    #30 c=1;//010->011 w=0->1 delay:132-120=12
    #30 c=0;//011->010 w=1->0 delay:162-150=12
    #30 a=1;//010->110 w=0->1 delay:199-180=19
    #30 b=0;//110->100 w=1->0 delay:227-210=17
    #30 c=1;//100->101 w=0->1 delay:252-240=12
    #30 c=0;//101->100 w=1->0 delay:282-270=12
    #30 b=1;//100->110 w=0->1 delay:319-300=19
    #30 a=0;//110->010 w=1->0 delay:347-330=17
    #30 $stop;
  end
endmodule